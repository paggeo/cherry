param int XLEN = 32;
param int OPSTART = 0;
param int OPSTOP = 6;
param int FUNCT3START = 12;
param int FUNCT3STOP = 14;
param int FUNCT7START = 25;
param int FUNCT7STOP = 31;

param int IMMSTART = 20;
param int IMMSTOP = 31;

param int SBFIRST_IMMSTART = 7;
param int SBFIRST_IMMSTOP = 11;
param int SBSECOND_IMMSTART = 25;
param int SBSECOND_IMMSTOP = 30;

param int UJFIRST_IMMSTART = 12;
param int UJFIRST_IMMSTOP = 19;

param int RDSTART = 7;
param int RDSTOP = 11;

param int RS1START = 15;
param int RS1STOP = 19;
param int RS2START = 20;
param int RS2STOP = 24;